module TC0030CMD(

);



endmodule
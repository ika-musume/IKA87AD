//this file defines microcode routine entrance

localparam NOP = 8'd255;